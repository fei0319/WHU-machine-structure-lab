module dm (
    input clk,
    input DMWr,
    input [5:0] address,
    input [31:0] din,
    input [2:0] DMType,
    output reg [31:0] dout
);

endmodule
